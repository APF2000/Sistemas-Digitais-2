library ieee;
use ieee.numeric_bit.all;

entity reg_tb is
end reg_tb;

architecture arc of reg_tb is

  flipFlop: process(clock, reset)
  begin

end arc;
